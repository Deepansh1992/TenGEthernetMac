package Macpackage
	`include *_sequence_item.sv
	`include *_sequence.sv
	`include *_driver.sv
	`include *_agent.sv
	`include monitor.sv
	`include environment.sv
endpackage