package pck; 
    `include *_sequence_item.sv
    `include *_sequence.sv
    `include *_driver.sv
    `include *_monitor.sv
    `include *_agent.sv
    // `include scoreboard.sv
    `include environment.sv
    `include testclass.sv
endpackage
    