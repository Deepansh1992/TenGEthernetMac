<<<<<<< HEAD
package pck; 
    `include *_sequence_item.sv
    `include *_sequence.sv
    `include *_driver.sv
    `include *_monitor.sv
    `include *_agent.sv
    // `include scoreboard.sv
    `include environment.sv
    `include testclass.sv
endpackage
    
=======
package Macpackage
	`include *_sequence_item.sv
	`include *_sequence.sv
	`include *_driver.sv
	`include *_agent.sv
	`include monitor.sv
	`include environment.sv
endpackage
>>>>>>> 80672db5b19edcfcb0382a5c07c37fa926f1ecb7
